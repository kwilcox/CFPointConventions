netcdf trajectoryProfile-Ragged-MultipleTrajectories-H.6.3 {
dimensions:
	obs = UNLIMITED ; // (548 currently)
	profile = 20 ;
	trajectory = 5 ;
variables:
	int trajectory(trajectory) ;
		trajectory:cf_role = "trajectory_id" ;
	float lat(profile) ;
		lat:units = "degrees_north" ;
		lat:long_name = "station latitude" ;
		lat:standard_name = "latitude" ;
	float lon(profile) ;
		lon:units = "degrees_east" ;
		lon:long_name = "station longitude" ;
		lon:standard_name = "longitude" ;
	int rowSize(profile) ;
		rowSize:long_name = "number of obs for this trajectory" ;
		rowSize:sample_dimension = "obs" ;
	int trajectory_index(profile) ;
		trajectory_index:long_name = "which trajectory this profile is for" ;
		trajectory_index:instance_dimension = "trajectory" ;
	int time(profile) ;
		time:long_name = "time of measurement" ;
		time:standard_name = "time" ;
		time:units = "seconds since 1990-01-01 00:00:00" ;
		time:missing_value = -999 ;
	float z(obs) ;
		z:long_name = "height above mean sea level" ;
		z:standard_name = "altitude" ;
		z:units = "m" ;
		z:positive = "up" ;
		z:axis = "Z" ;
		z:missing_value = -999.f ;
	float temperature(obs) ;
		temperature:long_name = "Air Temperature" ;
		temperature:standard_name = "air_temperature" ;
		temperature:units = "Celsius" ;
		temperature:coordinates = "time lat lon z" ;
		temperature:missing_value = -999.9f ;
	float humidity(obs) ;
		humidity:long_name = "Humidity" ;
		humidity:standard_name = "specific_humidity" ;
		humidity:units = "Percent" ;
		humidity:coordinates = "time lat lon z" ;
		humidity:missing_value = -999.9f ;

// global attributes:
		:Conventions = "CF-1.6" ;
		:featureType = "trajectoryProfile" ;
}
